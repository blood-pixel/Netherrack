module network

pub struct Network {

}

pub fn (mut n Network) init() {
    println("Network is starting")
}