module player