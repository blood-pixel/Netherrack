module world