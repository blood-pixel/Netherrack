module main

pub struct Netherrack {
}

pub fn (mut n Netherrack) start() {
}

fn main() {
    mut server := Netherrack{}
    server.start()
}