module entity